module u;
	always #1 $write("u");
endmodule